
-- Version-history: 

library ieee;
use ieee.std_logic_1164.all;

use work.lhc_data_pkg.all;
use work.gtl_pkg.all;

entity bx_pipeline is
    port(
        clk : in std_logic;
        data : in gtl_data_record;
        pt_muon_bx_p2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_muon_bx_p2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_muon_bx_p2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_muon_bx_p2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        qual_muon_bx_p2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        charge_muon_bx_p2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_muon_bx_p1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_muon_bx_p1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_muon_bx_p1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_muon_bx_p1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        qual_muon_bx_p1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        charge_muon_bx_p1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_muon_bx_0 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_muon_bx_0 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_muon_bx_0 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_muon_bx_0 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        qual_muon_bx_0 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        charge_muon_bx_0 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_muon_bx_m1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_muon_bx_m1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_muon_bx_m1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_muon_bx_m1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        qual_muon_bx_m1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        charge_muon_bx_m1 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_muon_bx_m2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_muon_bx_m2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_muon_bx_m2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_muon_bx_m2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        qual_muon_bx_m2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        charge_muon_bx_m2 : out obj_parameter_array(0 to MUON_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_eg_bx_p2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_eg_bx_p2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_eg_bx_p2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_eg_bx_p2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_eg_bx_p1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_eg_bx_p1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_eg_bx_p1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_eg_bx_p1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_eg_bx_0 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_eg_bx_0 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_eg_bx_0 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_eg_bx_0 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_eg_bx_m1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_eg_bx_m1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_eg_bx_m1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_eg_bx_m1 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_eg_bx_m2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_eg_bx_m2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_eg_bx_m2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_eg_bx_m2 : out obj_parameter_array(0 to EG_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_jet_bx_p2 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_jet_bx_p2 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_jet_bx_p2 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_jet_bx_p1 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_jet_bx_p1 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_jet_bx_p1 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_jet_bx_0 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_jet_bx_0 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_jet_bx_0 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_jet_bx_m1 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_jet_bx_m1 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_jet_bx_m1 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_jet_bx_m2 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_jet_bx_m2 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_jet_bx_m2 : out obj_parameter_array(0 to JET_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_tau_bx_p2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_tau_bx_p2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_tau_bx_p2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_tau_bx_p2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_tau_bx_p1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_tau_bx_p1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_tau_bx_p1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_tau_bx_p1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_tau_bx_0 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_tau_bx_0 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_tau_bx_0 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_tau_bx_0 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_tau_bx_m1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_tau_bx_m1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_tau_bx_m1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_tau_bx_m1 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        pt_tau_bx_m2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        eta_tau_bx_m2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        phi_tau_bx_m2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        iso_tau_bx_m2 : out obj_parameter_array(0 to TAU_ARRAY_LENGTH-1) := (others => (others => '0'));
        ett_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ett_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ett_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ett_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ett_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ht_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ht_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ht_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ht_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ht_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etm_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etm_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etm_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etm_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etm_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htm_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htm_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htm_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htm_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htm_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfp_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfp_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfp_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfp_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfp_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfm_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfm_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfm_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfm_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt1hfm_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfp_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfp_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfp_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfp_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfp_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfm_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfm_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfm_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfm_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        mbt0hfm_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ettem_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ettem_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ettem_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ettem_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        ettem_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etmhf_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etmhf_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etmhf_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etmhf_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        etmhf_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htmhf_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htmhf_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htmhf_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htmhf_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        htmhf_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        towercount_bx_p2 : out std_logic_vector(MAX_TOWERCOUNT_BITS-1 downto 0) := (others => '0');
        towercount_bx_p1 : out std_logic_vector(MAX_TOWERCOUNT_BITS-1 downto 0) := (others => '0');
        towercount_bx_0 : out std_logic_vector(MAX_TOWERCOUNT_BITS-1 downto 0) := (others => '0');
        towercount_bx_m1 : out std_logic_vector(MAX_TOWERCOUNT_BITS-1 downto 0) := (others => '0');
        towercount_bx_m2 : out std_logic_vector(MAX_TOWERCOUNT_BITS-1 downto 0) := (others => '0');
        asymet_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymet_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymet_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymet_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymet_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymht_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymht_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymht_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymht_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymht_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymethf_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymethf_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymethf_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymethf_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymethf_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymhthf_bx_p2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymhthf_bx_p1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymhthf_bx_0 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymhthf_bx_m1 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        asymhthf_bx_m2 : out std_logic_vector(MAX_ESUMS_BITS-1 downto 0) := (others => '0');
        centrality_bx_p2 : out std_logic_vector(NR_CENTRALITY_BITS-1 downto 0) := (others => '0');
        centrality_bx_p1 : out std_logic_vector(NR_CENTRALITY_BITS-1 downto 0) := (others => '0');
        centrality_bx_0 : out std_logic_vector(NR_CENTRALITY_BITS-1 downto 0) := (others => '0');
        centrality_bx_m1 : out std_logic_vector(NR_CENTRALITY_BITS-1 downto 0) := (others => '0');
        centrality_bx_m2 : out std_logic_vector(NR_CENTRALITY_BITS-1 downto 0) := (others => '0');
        ext_cond_bx_p2 : out std_logic_vector(EXTERNAL_CONDITIONS_DATA_WIDTH-1 downto 0) := (others => '0');
        ext_cond_bx_p1 : out std_logic_vector(EXTERNAL_CONDITIONS_DATA_WIDTH-1 downto 0) := (others => '0');
        ext_cond_bx_0 : out std_logic_vector(EXTERNAL_CONDITIONS_DATA_WIDTH-1 downto 0) := (others => '0');
        ext_cond_bx_m1 : out std_logic_vector(EXTERNAL_CONDITIONS_DATA_WIDTH-1 downto 0) := (others => '0');
        ext_cond_bx_m2 : out std_logic_vector(EXTERNAL_CONDITIONS_DATA_WIDTH-1 downto 0) := (others => '0')
    );
end bx_pipeline;

architecture rtl of bx_pipeline is

    constant pipeline_stages : natural := 5;
    type arr_eg_record_array is array (0 to pipeline_stages-1) of eg_record_array(0 to EG_ARRAY_LENGTH-1);    
    signal eg_bx_tmp : arr_eg_record_array;
    type arr_jet_record_array is array (0 to pipeline_stages-1) of jet_record_array(0 to JET_ARRAY_LENGTH-1);    
    signal jet_bx_tmp : arr_jet_record_array;
    type arr_tau_record_array is array (0 to pipeline_stages-1) of tau_record_array(0 to TAU_ARRAY_LENGTH-1);    
    signal tau_bx_tmp : arr_tau_record_array;
    type arr_muon_record_array is array (0 to pipeline_stages-1) of muon_record_array(0 to MUON_ARRAY_LENGTH-1);    
    signal muon_bx_tmp : arr_muon_record_array;

begin

    process(clk, data.eg_data, data.jet_data, data.tau_data, data.muon_data)
    begin
        eg_bx_tmp(0) <= data.eg_data;
        jet_bx_tmp(0) <= data.jet_data;
        tau_bx_tmp(0) <= data.tau_data;
        muon_bx_tmp(0) <= data.muon_data;
        for i in 0 to pipeline_stages-1-1 loop
            if (clk'event and clk = '1') then
                eg_bx_tmp(i+1) <= eg_bx_tmp(i);
                jet_bx_tmp(i+1) <= jet_bx_tmp(i);
                tau_bx_tmp(i+1) <= tau_bx_tmp(i);
                muon_bx_tmp(i+1) <= muon_bx_tmp(i);
            end if;
        end loop;
    end process;

    eg_l: for i in 0 to EG_ARRAY_LENGTH-1 generate
        pt_eg_bx_p2(i)(data.eg_data(i).pt'length-1 downto 0) <= eg_bx_tmp(0)(i).pt;
        eta_eg_bx_p2(i)(data.eg_data(i).eta'length-1 downto 0) <= eg_bx_tmp(0)(i).eta;
        phi_eg_bx_p2(i)(data.eg_data(i).phi'length-1 downto 0) <= eg_bx_tmp(0)(i).phi;
        iso_eg_bx_p2(i)(data.eg_data(i).iso'length-1 downto 0) <= eg_bx_tmp(0)(i).iso;
        pt_eg_bx_p1(i)(data.eg_data(i).pt'length-1 downto 0) <= eg_bx_tmp(1)(i).pt;
        eta_eg_bx_p1(i)(data.eg_data(i).eta'length-1 downto 0) <= eg_bx_tmp(1)(i).eta;
        phi_eg_bx_p1(i)(data.eg_data(i).phi'length-1 downto 0) <= eg_bx_tmp(1)(i).phi;
        iso_eg_bx_p1(i)(data.eg_data(i).iso'length-1 downto 0) <= eg_bx_tmp(1)(i).iso;
        pt_eg_bx_0(i)(data.eg_data(i).pt'length-1 downto 0) <= eg_bx_tmp(2)(i).pt;
        eta_eg_bx_0(i)(data.eg_data(i).eta'length-1 downto 0) <= eg_bx_tmp(2)(i).eta;
        phi_eg_bx_0(i)(data.eg_data(i).phi'length-1 downto 0) <= eg_bx_tmp(2)(i).phi;
        iso_eg_bx_0(i)(data.eg_data(i).iso'length-1 downto 0) <= eg_bx_tmp(2)(i).iso;
        pt_eg_bx_m1(i)(data.eg_data(i).pt'length-1 downto 0) <= eg_bx_tmp(3)(i).pt;
        eta_eg_bx_m1(i)(data.eg_data(i).eta'length-1 downto 0) <= eg_bx_tmp(3)(i).eta;
        phi_eg_bx_m1(i)(data.eg_data(i).phi'length-1 downto 0) <= eg_bx_tmp(3)(i).phi;
        iso_eg_bx_m1(i)(data.eg_data(i).iso'length-1 downto 0) <= eg_bx_tmp(3)(i).iso;
        pt_eg_bx_m2(i)(data.eg_data(i).pt'length-1 downto 0) <= eg_bx_tmp(4)(i).pt;
        eta_eg_bx_m2(i)(data.eg_data(i).eta'length-1 downto 0) <= eg_bx_tmp(4)(i).eta;
        phi_eg_bx_m2(i)(data.eg_data(i).phi'length-1 downto 0) <= eg_bx_tmp(4)(i).phi;
        iso_eg_bx_m2(i)(data.eg_data(i).iso'length-1 downto 0) <= eg_bx_tmp(4)(i).iso;
    end generate eg_l;

    jet_l: for i in 0 to JET_ARRAY_LENGTH-1 generate
        pt_jet_bx_p2(i)(data.jet_data(i).pt'length-1 downto 0) <= jet_bx_tmp(0)(i).pt;
        eta_jet_bx_p2(i)(data.jet_data(i).eta'length-1 downto 0) <= jet_bx_tmp(0)(i).eta;
        phi_jet_bx_p2(i)(data.jet_data(i).phi'length-1 downto 0) <= jet_bx_tmp(0)(i).phi;
        pt_jet_bx_p1(i)(data.jet_data(i).pt'length-1 downto 0) <= jet_bx_tmp(1)(i).pt;
        eta_jet_bx_p1(i)(data.jet_data(i).eta'length-1 downto 0) <= jet_bx_tmp(1)(i).eta;
        phi_jet_bx_p1(i)(data.jet_data(i).phi'length-1 downto 0) <= jet_bx_tmp(1)(i).phi;
        pt_jet_bx_0(i)(data.jet_data(i).pt'length-1 downto 0) <= jet_bx_tmp(2)(i).pt;
        eta_jet_bx_0(i)(data.jet_data(i).eta'length-1 downto 0) <= jet_bx_tmp(2)(i).eta;
        phi_jet_bx_0(i)(data.jet_data(i).phi'length-1 downto 0) <= jet_bx_tmp(2)(i).phi;
        pt_jet_bx_m1(i)(data.jet_data(i).pt'length-1 downto 0) <= jet_bx_tmp(3)(i).pt;
        eta_jet_bx_m1(i)(data.jet_data(i).eta'length-1 downto 0) <= jet_bx_tmp(3)(i).eta;
        phi_jet_bx_m1(i)(data.jet_data(i).phi'length-1 downto 0) <= jet_bx_tmp(3)(i).phi;
        pt_jet_bx_m2(i)(data.jet_data(i).pt'length-1 downto 0) <= jet_bx_tmp(4)(i).pt;
        eta_jet_bx_m2(i)(data.jet_data(i).eta'length-1 downto 0) <= jet_bx_tmp(4)(i).eta;
        phi_jet_bx_m2(i)(data.jet_data(i).phi'length-1 downto 0) <= jet_bx_tmp(4)(i).phi;
    end generate jet_l;

    tau_l: for i in 0 to TAU_ARRAY_LENGTH-1 generate
        pt_tau_bx_p2(i)(data.tau_data(i).pt'length-1 downto 0) <= tau_bx_tmp(0)(i).pt;
        eta_tau_bx_p2(i)(data.tau_data(i).eta'length-1 downto 0) <= tau_bx_tmp(0)(i).eta;
        phi_tau_bx_p2(i)(data.tau_data(i).phi'length-1 downto 0) <= tau_bx_tmp(0)(i).phi;
        iso_tau_bx_p2(i)(data.tau_data(i).iso'length-1 downto 0) <= tau_bx_tmp(0)(i).iso;
        pt_tau_bx_p1(i)(data.tau_data(i).pt'length-1 downto 0) <= tau_bx_tmp(1)(i).pt;
        eta_tau_bx_p1(i)(data.tau_data(i).eta'length-1 downto 0) <= tau_bx_tmp(1)(i).eta;
        phi_tau_bx_p1(i)(data.tau_data(i).phi'length-1 downto 0) <= tau_bx_tmp(1)(i).phi;
        iso_tau_bx_p1(i)(data.tau_data(i).iso'length-1 downto 0) <= tau_bx_tmp(1)(i).iso;
        pt_tau_bx_0(i)(data.tau_data(i).pt'length-1 downto 0) <= tau_bx_tmp(2)(i).pt;
        eta_tau_bx_0(i)(data.tau_data(i).eta'length-1 downto 0) <= tau_bx_tmp(2)(i).eta;
        phi_tau_bx_0(i)(data.tau_data(i).phi'length-1 downto 0) <= tau_bx_tmp(2)(i).phi;
        iso_tau_bx_0(i)(data.tau_data(i).iso'length-1 downto 0) <= tau_bx_tmp(2)(i).iso;
        pt_tau_bx_m1(i)(data.tau_data(i).pt'length-1 downto 0) <= tau_bx_tmp(3)(i).pt;
        eta_tau_bx_m1(i)(data.tau_data(i).eta'length-1 downto 0) <= tau_bx_tmp(3)(i).eta;
        phi_tau_bx_m1(i)(data.tau_data(i).phi'length-1 downto 0) <= tau_bx_tmp(3)(i).phi;
        iso_tau_bx_m1(i)(data.tau_data(i).iso'length-1 downto 0) <= tau_bx_tmp(3)(i).iso;
        pt_tau_bx_m2(i)(data.tau_data(i).pt'length-1 downto 0) <= tau_bx_tmp(4)(i).pt;
        eta_tau_bx_m2(i)(data.tau_data(i).eta'length-1 downto 0) <= tau_bx_tmp(4)(i).eta;
        phi_tau_bx_m2(i)(data.tau_data(i).phi'length-1 downto 0) <= tau_bx_tmp(4)(i).phi;
        iso_tau_bx_m2(i)(data.tau_data(i).iso'length-1 downto 0) <= tau_bx_tmp(4)(i).iso;
    end generate tau_l;

    muon_l: for i in 0 to MUON_ARRAY_LENGTH-1 generate
        pt_muon_bx_p2(i)(data.muon_data(i).pt'length-1 downto 0) <= muon_bx_tmp(0)(i).pt;
        eta_muon_bx_p2(i)(data.muon_data(i).eta'length-1 downto 0) <= muon_bx_tmp(0)(i).eta;
        phi_muon_bx_p2(i)(data.muon_data(i).phi'length-1 downto 0) <= muon_bx_tmp(0)(i).phi;
        iso_muon_bx_p2(i)(data.muon_data(i).iso'length-1 downto 0) <= muon_bx_tmp(0)(i).iso;
        qual_muon_bx_p2(i)(data.muon_data(i).qual'length-1 downto 0) <= muon_bx_tmp(0)(i).qual;
        charge_muon_bx_p2(i)(data.muon_data(i).charge'length-1 downto 0) <= muon_bx_tmp(0)(i).charge;
        pt_muon_bx_p1(i)(data.muon_data(i).pt'length-1 downto 0) <= muon_bx_tmp(1)(i).pt;
        eta_muon_bx_p1(i)(data.muon_data(i).eta'length-1 downto 0) <= muon_bx_tmp(1)(i).eta;
        phi_muon_bx_p1(i)(data.muon_data(i).phi'length-1 downto 0) <= muon_bx_tmp(1)(i).phi;
        iso_muon_bx_p1(i)(data.muon_data(i).iso'length-1 downto 0) <= muon_bx_tmp(1)(i).iso;
        qual_muon_bx_p1(i)(data.muon_data(i).qual'length-1 downto 0) <= muon_bx_tmp(1)(i).qual;
        charge_muon_bx_p1(i)(data.muon_data(i).charge'length-1 downto 0) <= muon_bx_tmp(1)(i).charge;
        pt_muon_bx_0(i)(data.muon_data(i).pt'length-1 downto 0) <= muon_bx_tmp(2)(i).pt;
        eta_muon_bx_0(i)(data.muon_data(i).eta'length-1 downto 0) <= muon_bx_tmp(2)(i).eta;
        phi_muon_bx_0(i)(data.muon_data(i).phi'length-1 downto 0) <= muon_bx_tmp(2)(i).phi;
        iso_muon_bx_0(i)(data.muon_data(i).iso'length-1 downto 0) <= muon_bx_tmp(2)(i).iso;
        qual_muon_bx_0(i)(data.muon_data(i).qual'length-1 downto 0) <= muon_bx_tmp(2)(i).qual;
        charge_muon_bx_0(i)(data.muon_data(i).charge'length-1 downto 0) <= muon_bx_tmp(2)(i).charge;
        pt_muon_bx_m1(i)(data.muon_data(i).pt'length-1 downto 0) <= muon_bx_tmp(3)(i).pt;
        eta_muon_bx_m1(i)(data.muon_data(i).eta'length-1 downto 0) <= muon_bx_tmp(3)(i).eta;
        phi_muon_bx_m1(i)(data.muon_data(i).phi'length-1 downto 0) <= muon_bx_tmp(3)(i).phi;
        iso_muon_bx_m1(i)(data.muon_data(i).iso'length-1 downto 0) <= muon_bx_tmp(3)(i).iso;
        qual_muon_bx_m1(i)(data.muon_data(i).qual'length-1 downto 0) <= muon_bx_tmp(3)(i).qual;
        charge_muon_bx_m1(i)(data.muon_data(i).charge'length-1 downto 0) <= muon_bx_tmp(3)(i).charge;
        pt_muon_bx_m2(i)(data.muon_data(i).pt'length-1 downto 0) <= muon_bx_tmp(4)(i).pt;
        eta_muon_bx_m2(i)(data.muon_data(i).eta'length-1 downto 0) <= muon_bx_tmp(4)(i).eta;
        phi_muon_bx_m2(i)(data.muon_data(i).phi'length-1 downto 0) <= muon_bx_tmp(4)(i).phi;
        iso_muon_bx_m2(i)(data.muon_data(i).iso'length-1 downto 0) <= muon_bx_tmp(4)(i).iso;
        qual_muon_bx_m2(i)(data.muon_data(i).qual'length-1 downto 0) <= muon_bx_tmp(4)(i).qual;
        charge_muon_bx_m2(i)(data.muon_data(i).charge'length-1 downto 0) <= muon_bx_tmp(4)(i).charge;
    end generate muon_l;

end architecture rtl;
